`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:39:23 08/26/2015 
// Design Name: 
// Module Name:    Sincronizador 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

	/* 
	 *Modulo encargado de sincronizar las entradas con el reloj del sistema.
	 *Tiene como entradas 3 bits del identificador del piso en código Gray, la señal
	 *binaria del sensor de sobrepeso, la señal binaria del sensor de obtaculización de la puerta
	 *y los 2 bits por cada uno de los 5 pisos donde el MSB es señal desubida y el LSB de bajada
	 */
	 
module Sincronizador(
    );


endmodule
