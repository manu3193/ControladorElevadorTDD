`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:33:57 08/26/2015 
// Design Name: 
// Module Name:    DivisorFrecuencia 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////


  /*
	*Este módulo recibe como entrada el clock del dispositivo e implementa un divisor de
	*de frecuencias con sumadores binarios que da como salida el reloj del sistema
	*controlador del ascensor, a 1 Hz. 
	*
   */

module DivisorFrecuencia(
    );


endmodule
