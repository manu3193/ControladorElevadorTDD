`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:31:03 08/26/2015 
// Design Name: 
// Module Name:    RegistroSolicitudes 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////


	/*
	 *Este módulo se encarga de registrar las solucitudes de todos los pisos
	 *implementando un banco de 5 registros de 2 bits secuenciales, activados 
	 *por un mismo reloj.
	 *Tiene como entrada 5 pares de 2 bits.
	 *
	 */
module RegistroSolicitudes(
    );


endmodule
