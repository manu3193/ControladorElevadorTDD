`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:33:33 08/26/2015 
// Design Name: 
// Module Name:    VerificadorSentidoMovimiento 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////


	/*
	 *Módulo encargado de decidir el movimiendo y la dirección del ascensor mediante
	 *lógica combinacional entre el valor del registro de solicitudes y el piso actual.
	 *Tiene como entradas los 10 bits del registro de solicitudes y los 3 bits del código
	 *Grey identificador de cada piso y el clock. Tiene como salidas 2 bits que idicarán la
	 *habilitación del motor (MSB) 0=apagado, 1=activado y la dirección(LSB) 0=bajar, 1=subir . 
	 */
	 
module VerificadorSentidoMovimiento(
    );


endmodule
