`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   23:37:41 08/26/2015
// Design Name:   DecoBCDto7seg
// Module Name:   /home/manzumbado/Development/HDL/Xilinx/ControladorElevadorTDD/trunk/DecoGreytoBCD.v
// Project Name:  ControladorElevadorTDD
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: DecoBCDto7seg
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module DecoGreytoBCD;

      
endmodule

