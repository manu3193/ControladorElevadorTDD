`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:33:03 08/26/2015 
// Design Name: 
// Module Name:    Temporizador 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

	/*
	 *Módulo encargado de implementar un temporizador. Tiene como entradas una señal de inicio,
	 *una señal de restart y la entrada de reloj del sistema. Como salida debe retornar una señal 
	 *que se active cuando termina de contar el tiempo definido.
	 *
	 */
	 
module Temporizador(
    );


endmodule
